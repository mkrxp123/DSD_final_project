`include "CONSTANT.v"

// module matrix_mul #(parameter WIDTH = `MAX_WIDTH) (
//     input
// );
    
// endmodule