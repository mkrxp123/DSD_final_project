`include "element_op.v"

module tb ();

endmodule