`include "CONSTANT.v"
`include "processor.v"

module tb ();
    
endmodule